----------------------------------------------------------------------------------
-- Name:	Prof Jeff Falkinburg
-- Date:	Fall 2020
-- Course:	CSCE 230
-- File:	SimpleComputer.vhd
-- HW:		Group Project
-- Purp:	Implements the top-level design of our Simple Computer for our project 
--
-- Doc:		Lecture Notes
-- 	
-- Academic Integrity Statement: I certify that, while others may have 
-- assisted me in brain storming, debugging and validating this program, 
-- the program itself is my own work. I understand that submitting code 
-- which is the work of other individuals is a violation of the honor   
-- code.  I also understand that if I knowingly give my original work to 
-- another individual is also a violation of the honor code. 
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

entity SimpleComputer is
	port(
		clock			: in std_logic;
		LEDR 			: out std_logic_vector(9 downto 0);
		HEX_DP		: out std_logic_vector(7 downto 0);
		SW 			: in std_logic_vector(9 downto 0);
		KEY 			: in std_logic_vector(1 downto 0):= "10"; -- reset = not KEY0
		-- for ModelSim debugging only
		debug_PC	: out std_logic_vector(15 downto 0);
		debug_IR	: out std_logic_vector(15 downto 0);
		debug_state : out std_logic_vector(2 downto 0);
		debug_r1	: out std_logic_vector(15 downto 0);
		debug_r2	: out std_logic_vector(15 downto 0);
		debug_r3	: out std_logic_vector(15 downto 0);
		debug_r4	: out std_logic_vector(15 downto 0);
		debug_r5	: out std_logic_vector(15 downto 0);
		debug_r6	: out std_logic_vector(15 downto 0);
		debug_r7	: out std_logic_vector(15 downto 0);
		debug_RA	: out std_logic_vector(15 downto 0);
		debug_RB	: out std_logic_vector(15 downto 0);
		debug_Extension : out std_logic_vector(15 downto 0);
		debug_RZ	: out std_logic_vector(15 downto 0);
		debug_RY	: out std_logic_vector(15 downto 0)
	);
end SimpleComputer;

architecture implementation of SimpleComputer is
	component SimpleProcessor is
		port(
			clock			: in std_logic;
			reset			: in std_logic;
			MEM_read		: out std_logic;
			MEM_write	: out std_logic;
			MFC			: in std_logic;
			MEM_address	: out std_logic_vector(15 downto 0);
			Data_to_Mem	: out std_logic_vector(15 downto 0);
			Data_from_Mem : in std_logic_vector(15 downto 0);
			-- for ModelSim debugging only
			debug_PC	: out std_logic_vector(15 downto 0);
			debug_IR	: out std_logic_vector(15 downto 0);
			debug_state : out std_logic_vector(2 downto 0);
			debug_r1	: out std_logic_vector(15 downto 0);
			debug_r2	: out std_logic_vector(15 downto 0);
			debug_r3	: out std_logic_vector(15 downto 0);
			debug_r4	: out std_logic_vector(15 downto 0);
			debug_r5	: out std_logic_vector(15 downto 0);
			debug_r6	: out std_logic_vector(15 downto 0);
			debug_r7	: out std_logic_vector(15 downto 0);
			debug_RA	: out std_logic_vector(15 downto 0);
			debug_RB	: out std_logic_vector(15 downto 0);
			debug_Extension : out std_logic_vector(15 downto 0);
			debug_RZ	: out std_logic_vector(15 downto 0);
			debug_RY	: out std_logic_vector(15 downto 0);
			debug_adder	: out std_logic_vector(15 downto 0)
		);
	end component;
	component MemoryIOInterface is
		port(
			clock 		: in std_logic;
			reset			: in std_logic;
			MEM_read		: in std_logic;
			MEM_write 	: in std_logic;
			MFC			: out std_logic;
			Address 		: in std_logic_vector(15 downto 0);
			Data_in 		: in std_logic_vector(15 downto 0);
			Data_out		: out std_logic_vector(15 downto 0);
			LEDR 			: out std_logic_vector(9 downto 0);
			HEX_DP 		: out std_logic_vector(7 downto 0);
			SW 			: in std_logic_vector(9 downto 0);
			KEY 			: in std_logic
		);
	end component;
	
	signal	MFC, MEM_read, MEM_write: std_logic;
	signal	Address, Data_from_Mem, Data_to_Mem: std_logic_vector(15 downto 0);
	signal	debug_adder : std_logic_vector(15 downto 0);
begin

	-- processor uses the rising edge, and is reset when pushing KEY0
	P: SimpleProcessor port map (clock=>clock, reset=>not KEY(0), 
			MEM_read=>MEM_read, MEM_write=>MEM_write,
			MFC=>MFC, MEM_address=>Address,
			Data_to_Mem=>Data_to_Mem, Data_from_Mem=>Data_from_Mem,
			debug_PC=>debug_PC, debug_IR=>debug_IR, debug_state=>debug_state,
			debug_r1=>debug_r1, debug_r2=>debug_r2, debug_r3=>debug_r3,
			debug_r4=>debug_r4, debug_r5=>debug_r5, debug_r6=>debug_r6, debug_r7=>debug_r7,
			debug_RA=>debug_RA, debug_RB=>debug_RB, debug_Extension=>debug_Extension,
			debug_RZ=>debug_RZ, debug_RY=>debug_RY, debug_adder=>debug_adder);
					
	
	-- memory and IO use the falling edge, and is reset when pushing KEY0
	MemIO: MemoryIOInterface port map (clock=>not clock, reset=>not KEY(0), 
			MEM_read=>MEM_read, MEM_write=>MEM_write,
			MFC=>MFC, Address=>Address, 
			Data_in=>Data_to_Mem, Data_out=>Data_from_Mem,
			KEY=>KEY(1), SW=>SW, HEX_DP=>HEX_DP, LEDR=>LEDR);
			
end implementation;
